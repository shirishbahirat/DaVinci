/*
File Name   : Test_ALU.v
Description : RISC-V RV32I 算数逻辑单元 测试
Written By  : Tealer Guo
Data        : 2019/04/20
*/
`timescale 1ns/1ns
// 测试模块
module alu_test;
	reg[31:0] rs1_num;
	reg[31:0] rs2_num;
	// ALU操作数
	reg[9:0] alu_op;
	// 结果
	wire[31:0] rd_num;
	// 实例化模块
	ALU alu_test(
		.rs1_num(rs1_num),
		.rs2_num(rs2_num),
		.alu_op(alu_op),
		.rd_num(rd_num)
	);
	// 仿真设置
	// 32-bit 00000000000000000000000000000000
	initial
		begin
			#0 rs1_num=32'b00000000000010000010001010010110;rs2_num=32'b01000001111000010111100100110110;alu_op=10'b0000000001;//and
			#5 rs1_num=32'b01001100000010010010000100011010;rs2_num=32'b00000000001000010101100100110100;alu_op=10'b0000000010;//sub
			#5 rs1_num=32'b10000010010010010010100010011100;rs2_num=32'b00010001101001010000100000110010;alu_op=10'b0000001001;//sra
			#5 rs1_num=32'b00100010000010001010001000010110;rs2_num=32'b01010001011011111000100100110011;alu_op=10'b0000001010;//or
			#5 rs1_num=32'b00000100000010100010010010011000;rs2_num=32'b00110001001000010100100100111111;alu_op=10'b0000000001;//and
			#5 rs1_num=32'b00000000000010000010001010010110;rs2_num=32'b01000001111000010111100100110110;alu_op=10'b0000000011;//sll
			#5 rs1_num=32'b01001100000010010010000100011010;rs2_num=32'b00000000001000010101100100110100;alu_op=10'b0000000101;//slt
			#5 rs1_num=32'b00000010010010010010100010011100;rs2_num=32'b00010001101001010000100000110010;alu_op=10'b0000000110;//sltu
			#5 rs1_num=32'b00100010000010001010001000010110;rs2_num=32'b01010001011011111000100100110011;alu_op=10'b0000000111;//xor
			#5 rs1_num=32'b00000100000010100010010010011000;rs2_num=32'b00110001001000010100100100111111;alu_op=10'b0000001000;//srl
			#5 $finish;
		end
	// vvp设置
	initial
		begin
			$dumpfile("ALU.vcd");
			$dumpvars(0,alu_test);
		end

endmodule